.subckt an21 A B VDD VSS Y
M5 Y net26 VSS VSS NMOS w=2u l=1u
M4 N001 A VSS VSS NMOS w=2u l=1u
M3 net26 B N001 VSS NMOS w=2u l=1u
M2 Y net26 VDD VDD PMOS w=6u l=1u
M1 net26 B VDD VDD PMOS w=6u l=1u
M0 net26 A VDD VDD PMOS w=6u l=1u
.ends an21

.subckt an31 A B C VDD VSS Y
M7 Y net19 VDD VDD PMOS w=6u l=1u
M6 net19 C VDD VDD PMOS w=6u l=1u
M5 net19 B VDD VDD PMOS w=6u l=1u
M4 net19 A VDD VDD PMOS w=6u l=1u
M3 Y net19 VSS VSS NMOS w=2u l=1u
M2 net19 C N001 VSS NMOS w=4.7u l=1u
M1 N001 B N002 VSS NMOS w=4.7u l=1u
M0 N002 A VSS VSS NMOS w=4.7u l=1u
.ends an31

.subckt an41 A B C D VDD VSS Y
M8 Y net44 VSS VSS NMOS w=2u l=1u
M7 N003 A VSS VSS NMOS w=6.2u l=1u
M6 N002 B N003 VSS NMOS w=6.2u l=1u
M5 N001 C N002 VSS NMOS w=6.2u l=1u
M4 net44 D N001 VSS NMOS w=6.2u l=1u
M9 Y net44 VDD VDD PMOS w=6u l=1u
M3 net44 D VDD VDD PMOS w=6u l=1u
M2 net44 C VDD VDD PMOS w=6u l=1u
M1 net44 B VDD VDD PMOS w=6u l=1u
M0 net44 A VDD VDD PMOS w=6u l=1u
.ends an41

.subckt buf1 A VDD VSS Y
M3 Y net13 VDD VDD PMOS w=6u l=1u
M2 net13 A VDD VDD PMOS w=6u l=1u
M1 net13 A VSS VSS NMOS w=2u l=1u
M0 Y net13 VSS VSS NMOS w=2u l=1u
.ends buf1

.subckt buf2 A VDD VSS Y
M4 Y net13 VDD VDD PMOS w=6u l=1u
M3 Y net13 VDD VDD PMOS w=6u l=1u
M2 net13 A VDD VDD PMOS w=6u l=1u
M5 Y net13 VSS VSS NMOS w=2u l=1u
M1 net13 A VSS VSS NMOS w=2u l=1u
M0 Y net13 VSS VSS NMOS w=2u l=1u
.ends buf2

.subckt buf4 A VDD VSS Y
M8 Y net13 VDD VDD PMOS w=6u l=1u
M6 Y net13 VDD VDD PMOS w=6u l=1u
M4 Y net13 VDD VDD PMOS w=6u l=1u
M3 Y net13 VDD VDD PMOS w=6u l=1u
M2 net13 A VDD VDD PMOS w=6u l=1u
M9 Y net13 VSS VSS NMOS w=2u l=1u
M7 Y net13 VSS VSS NMOS w=2u l=1u
M5 Y net13 VSS VSS NMOS w=2u l=1u
M1 net13 A VSS VSS NMOS w=2u l=1u
M0 Y net13 VSS VSS NMOS w=2u l=1u
.ends buf4

.subckt buf8 A VDD VSS Y
M17 Y net13 VDD VDD PMOS w=6u l=1u
M15 Y net13 VDD VDD PMOS w=6u l=1u
M12 Y net13 VDD VDD PMOS w=6u l=1u
M10 Y net13 VDD VDD PMOS w=6u l=1u
M8 Y net13 VDD VDD PMOS w=6u l=1u
M6 Y net13 VDD VDD PMOS w=6u l=1u
M4 Y net13 VDD VDD PMOS w=6u l=1u
M3 Y net13 VDD VDD PMOS w=6u l=1u
M2 net13 A VDD VDD PMOS w=6u l=1u
M16 Y net13 VSS VSS NMOS w=2u l=1u
M14 Y net13 VSS VSS NMOS w=2u l=1u
M13 Y net13 VSS VSS NMOS w=2u l=1u
M11 Y net13 VSS VSS NMOS w=2u l=1u
M9 Y net13 VSS VSS NMOS w=2u l=1u
M7 Y net13 VSS VSS NMOS w=2u l=1u
M5 Y net13 VSS VSS NMOS w=2u l=1u
M1 net13 A VSS VSS NMOS w=2u l=1u
M0 Y net13 VSS VSS NMOS w=2u l=1u
.ends buf8

.subckt cinv A OE VDD VSS YB
M5 net6 OE VSS VSS NMOS w=2u l=1u
M4 N002 A VSS VSS NMOS w=2u l=1u
M3 YB OE N002 VSS NMOS w=2u l=1u
M2 net6 OE VDD VDD PMOS w=6u l=1u
M1 YB net6 N001 VDD PMOS w=6u l=1u
M0 N001 A VDD VDD PMOS w=6u l=1u
.ends cinv

.subckt clkbuf2 A VDD VSS Y
M4 Y net13 VDD VDD PMOS w=6u l=1u
M3 Y net13 VDD VDD PMOS w=6u l=1u
M2 net13 A VDD VDD PMOS w=6u l=1u
M5 Y net13 VSS VSS NMOS w=2.4u l=1u
M1 net13 A VSS VSS NMOS w=2.4u l=1u
M0 Y net13 VSS VSS NMOS w=2.4u l=1u
.ends clkbuf2

.subckt clkinv1 A VDD VSS YB
M3 YB A VDD VDD PMOS w=6u l=1u
M0 YB A VSS VSS NMOS w=2.4u l=1u
.ends clkinv1

.subckt clkinv2 A VDD VSS YB
M4 YB A VDD VDD PMOS w=6u l=1u
M3 YB A VDD VDD PMOS w=6u l=1u
M5 YB A VSS VSS NMOS w=2.4u l=1u
M0 YB A VSS VSS NMOS w=2.4u l=1u
.ends clkinv2

.subckt dff1 CK D Q VDD VSS
M26 Q net66 VDD VDD PMOS w=6u l=1u
M24 net66 net92 VDD VDD PMOS w=6u l=1u
M18 net78 net116 N003 VDD PMOS w=6u l=1u
M17 net78 net74 N004 VDD PMOS w=6u l=1u
M16 N003 net104 VDD VDD PMOS w=6u l=1u
M15 N004 net92 VDD VDD PMOS w=6u l=1u
M14 net92 net78 VDD VDD PMOS w=6u l=1u
M13 net104 net114 VDD VDD PMOS w=6u l=1u
M12 N002 net104 VDD VDD PMOS w=6u l=1u
M11 N001 D VDD VDD PMOS w=6u l=1u
M10 net114 net116 N002 VDD PMOS w=6u l=1u
M9 net114 net74 N001 VDD PMOS w=6u l=1u
M8 net116 net74 VDD VDD PMOS w=6u l=1u
M7 net74 CK VDD VDD PMOS w=6u l=1u
M27 Q net66 VSS VSS NMOS w=2u l=1u
M25 net66 net92 VSS VSS NMOS w=2u l=1u
M23 net78 net74 N007 VSS NMOS w=2u l=1u
M22 N007 net104 VSS VSS NMOS w=2u l=1u
M21 net78 net116 N008 VSS NMOS w=2u l=1u
M20 N008 net92 VSS VSS NMOS w=2u l=1u
M19 net92 net78 VSS VSS NMOS w=2u l=1u
M6 net116 net74 VSS VSS NMOS w=2u l=1u
M5 net74 CK VSS VSS NMOS w=2u l=1u
M4 net104 net114 VSS VSS NMOS w=2u l=1u
M3 N006 net104 VSS VSS NMOS w=2u l=1u
M2 net114 net74 N006 VSS NMOS w=2u l=1u
M1 N005 D VSS VSS NMOS w=2u l=1u
M0 net114 net116 N005 VSS NMOS w=2u l=1u
.ends dff1

.subckt exnr A B VDD VSS YB
M9 net18 B VSS VSS NMOS w=2u l=1u
M8 net18 A VSS VSS NMOS w=2u l=1u
M7 YB net42 net18 VSS NMOS w=2u l=1u
M6 N002 B VSS VSS NMOS w=2u l=1u
M5 net42 A N002 VSS NMOS w=2u l=1u
M4 YB net42 VDD VDD PMOS w=6u l=1u
M3 YB B N001 VDD PMOS w=6u l=1u
M2 N001 A VDD VDD PMOS w=6u l=1u
M1 net42 B VDD VDD PMOS w=6u l=1u
M0 net42 A VDD VDD PMOS w=6u l=1u
.ends exnr

.subckt exor A B VDD VSS Y
M9 net106 A VDD VDD PMOS w=6u l=1u
M8 net106 B VDD VDD PMOS w=6u l=1u
M7 Y net134 net106 VDD PMOS w=6u l=1u
M6 N001 A VDD VDD PMOS w=6u l=1u
M5 net134 B N001 VDD PMOS w=6u l=1u
M4 Y net134 VSS VSS NMOS w=2u l=1u
M3 N002 B VSS VSS NMOS w=2u l=1u
M2 Y A N002 VSS NMOS w=2u l=1u
M1 net134 B VSS VSS NMOS w=2u l=1u
M0 net134 A VSS VSS NMOS w=2u l=1u
.ends exor

.subckt inv1 A VDD VSS YB
M3 YB A VDD VDD PMOS w=6u l=1u
M0 YB A VSS VSS NMOS w=2u l=1u
.ends inv1

.subckt inv2 A VDD VSS YB
M4 YB A VDD VDD PMOS w=6u l=1u
M3 YB A VDD VDD PMOS w=6u l=1u
M5 YB A VSS VSS NMOS w=2u l=1u
M0 YB A VSS VSS NMOS w=2u l=1u
.ends inv2

.subckt inv4 A VDD VSS YB
M8 YB A VDD VDD PMOS w=6u l=1u
M6 YB A VDD VDD PMOS w=6u l=1u
M4 YB A VDD VDD PMOS w=6u l=1u
M3 YB A VDD VDD PMOS w=6u l=1u
M9 YB A VSS VSS NMOS w=2u l=1u
M7 YB A VSS VSS NMOS w=2u l=1u
M5 YB A VSS VSS NMOS w=2u l=1u
M0 YB A VSS VSS NMOS w=2u l=1u
.ends inv4

.subckt inv8 A VDD VSS YB
M17 YB A VDD VDD PMOS w=6u l=1u
M15 YB A VDD VDD PMOS w=6u l=1u
M12 YB A VDD VDD PMOS w=6u l=1u
M10 YB A VDD VDD PMOS w=6u l=1u
M8 YB A VDD VDD PMOS w=6u l=1u
M6 YB A VDD VDD PMOS w=6u l=1u
M4 YB A VDD VDD PMOS w=6u l=1u
M3 YB A VDD VDD PMOS w=6u l=1u
M16 YB A VSS VSS NMOS w=2u l=1u
M14 YB A VSS VSS NMOS w=2u l=1u
M13 YB A VSS VSS NMOS w=2u l=1u
M11 YB A VSS VSS NMOS w=2u l=1u
M9 YB A VSS VSS NMOS w=2u l=1u
M7 YB A VSS VSS NMOS w=2u l=1u
M5 YB A VSS VSS NMOS w=2u l=1u
M0 YB A VSS VSS NMOS w=2u l=1u
.ends inv8

.subckt na212 A0 A1 B0 VDD VSS YB
M5 net031 A1 VSS VSS NMOS w=2u l=1u
M4 net031 A0 VSS VSS NMOS w=2u l=1u
M3 YB B0 net031 VSS NMOS w=2u l=1u
M2 YB B0 VDD VDD PMOS w=6u l=1u
M1 YB A1 N001 VDD PMOS w=6u l=1u
M0 N001 A0 VDD VDD PMOS w=6u l=1u
.ends na212

.subckt na21 A B VDD VSS YB
M4 N001 A VSS VSS NMOS w=2u l=1u
M3 YB B N001 VSS NMOS w=2u l=1u
M1 YB B VDD VDD PMOS w=6u l=1u
M0 YB A VDD VDD PMOS w=6u l=1u
.ends na21

.subckt na222 A0 A1 B0 B1 VDD VSS YB
M7 net12 A1 VSS VSS NMOS w=2u l=1u
M6 net12 A0 VSS VSS NMOS w=2u l=1u
M5 YB B1 net12 VSS NMOS w=2u l=1u
M4 YB B0 net12 VSS NMOS w=2u l=1u
M3 YB A1 N002 VDD PMOS w=6u l=1u
M2 N002 A0 VDD VDD PMOS w=6u l=1u
M1 YB B1 N001 VDD PMOS w=6u l=1u
M0 N001 B0 VDD VDD PMOS w=6u l=1u
.ends na222

.subckt na31 A B C VDD VSS YB
M6 YB C VDD VDD PMOS w=6u l=1u
M5 YB B VDD VDD PMOS w=6u l=1u
M4 YB A VDD VDD PMOS w=6u l=1u
M2 YB C N001 VSS NMOS w=4.7u l=1u
M1 N001 B N002 VSS NMOS w=4.7u l=1u
M0 N002 A VSS VSS NMOS w=4.7u l=1u
.ends na31

.subckt na41 A B C D VDD VSS YB
M7 N003 A VSS VSS NMOS w=6.2u l=1u
M6 N002 B N003 VSS NMOS w=6.2u l=1u
M5 N001 C N002 VSS NMOS w=6.2u l=1u
M4 YB D N001 VSS NMOS w=6.2u l=1u
M3 YB D VDD VDD PMOS w=6u l=1u
M2 YB C VDD VDD PMOS w=6u l=1u
M1 YB B VDD VDD PMOS w=6u l=1u
M0 YB A VDD VDD PMOS w=6u l=1u
.ends na41

.subckt nr212 A0 A1 B0 VDD VSS YB
M5 net18 A1 VDD VDD PMOS w=6u l=1u
M4 net18 A0 VDD VDD PMOS w=6u l=1u
M3 YB B0 net18 VDD PMOS w=6u l=1u
M2 YB B0 VSS VSS NMOS w=2u l=1u
M1 N001 A0 VSS VSS NMOS w=2u l=1u
M0 YB A1 N001 VSS NMOS w=2u l=1u
.ends nr212

.subckt nr21 A B VDD VSS YB
M3 N001 A VDD VDD PMOS w=6u l=1u
M2 YB B N001 VDD PMOS w=6u l=1u
M1 YB B VSS VSS NMOS w=2u l=1u
M0 YB A VSS VSS NMOS w=2u l=1u
.ends nr21

.subckt nr222 A0 A1 B0 B1 VDD VSS YB
M7 N001 A0 VSS VSS NMOS w=2u l=1u
M6 N002 B0 VSS VSS NMOS w=2u l=1u
M5 YB B1 N002 VSS NMOS w=2u l=1u
M4 YB A1 N001 VSS NMOS w=2u l=1u
M3 YB B1 net31 VDD PMOS w=6u l=1u
M2 YB B0 net31 VDD PMOS w=6u l=1u
M1 net31 A1 VDD VDD PMOS w=6u l=1u
M0 net31 A0 VDD VDD PMOS w=6u l=1u
.ends nr222

.subckt nr31 A B C VDD VSS YB
M5 YB C VSS VSS NMOS w=2u l=1u
M4 YB B VSS VSS NMOS w=2u l=1u
M3 YB A VSS VSS NMOS w=2u l=1u
M2 YB C N002 VDD PMOS w=12.6u l=1u
M1 N002 B N001 VDD PMOS w=12.6u l=1u
M0 N001 A VDD VDD PMOS w=12.6u l=1u
.ends nr31

.subckt or21 A B VDD VSS Y
M4 Y net068 VDD VDD PMOS w=6u l=1u
M3 N001 A VDD VDD PMOS w=6u l=1u
M2 net068 B N001 VDD PMOS w=6u l=1u
M5 Y net068 VSS VSS NMOS w=2u l=1u
M1 net068 B VSS VSS NMOS w=2u l=1u
M0 net068 A VSS VSS NMOS w=2u l=1u
.ends or21

.subckt or31 A B C VDD VSS Y
M7 Y net075 VSS VSS NMOS w=2u l=1u
M5 net075 C VSS VSS NMOS w=2u l=1u
M4 net075 B VSS VSS NMOS w=2u l=1u
M3 net075 A VSS VSS NMOS w=2u l=1u
M6 Y net075 VDD VDD PMOS w=6u l=1u
M2 net075 C N002 VDD PMOS w=12.6u l=1u
M1 N002 B N001 VDD PMOS w=12.6u l=1u
M0 N001 A VDD VDD PMOS w=12.6u l=1u
.ends or31

.subckt rff1 CK D Q QB R VDD VSS
M29 net104 R N003 VDD PMOS w=6u l=1u
M31 net92 R N006 VDD PMOS w=6u l=1u
M26 Q QB VDD VDD PMOS w=6u l=1u
M24 QB net92 VDD VDD PMOS w=6u l=1u
M18 net78 net116 N004 VDD PMOS w=6u l=1u
M17 net78 net74 N005 VDD PMOS w=6u l=1u
M16 N004 net104 VDD VDD PMOS w=6u l=1u
M15 N005 net92 VDD VDD PMOS w=6u l=1u
M14 N006 net78 VDD VDD PMOS w=6u l=1u
M13 N003 net114 VDD VDD PMOS w=6u l=1u
M12 N002 net104 VDD VDD PMOS w=6u l=1u
M11 N001 D VDD VDD PMOS w=6u l=1u
M10 net114 net116 N002 VDD PMOS w=6u l=1u
M9 net114 net74 N001 VDD PMOS w=6u l=1u
M8 net116 net74 VDD VDD PMOS w=6u l=1u
M7 net74 CK VDD VDD PMOS w=6u l=1u
M27 Q QB VSS VSS NMOS w=2u l=1u
M25 QB net92 VSS VSS NMOS w=2u l=1u
M23 net78 net74 N009 VSS NMOS w=2u l=1u
M22 N009 net104 VSS VSS NMOS w=2u l=1u
M21 net78 net116 N010 VSS NMOS w=2u l=1u
M20 N010 net92 VSS VSS NMOS w=2u l=1u
M19 net92 net78 VSS VSS NMOS w=2u l=1u
M30 net92 R VSS VSS NMOS w=2u l=1u
M28 net104 R VSS VSS NMOS w=2u l=1u
M6 net116 net74 VSS VSS NMOS w=2u l=1u
M5 net74 CK VSS VSS NMOS w=2u l=1u
M4 net104 net114 VSS VSS NMOS w=2u l=1u
M3 N008 net104 VSS VSS NMOS w=2u l=1u
M2 net114 net74 N008 VSS NMOS w=2u l=1u
M1 N007 D VSS VSS NMOS w=2u l=1u
M0 net114 net116 N007 VSS NMOS w=2u l=1u
.ends rff1

.subckt sdff1 CK D Q SE SI VDD VSS
M39 net0275 net0287 VDD VDD PMOS w=6u l=1u
M28 net0367 SE VDD VDD PMOS w=6u l=1u
M32 net0287 D VDD VDD PMOS w=6u l=1u
M33 net0287 net0367 VDD VDD PMOS w=6u l=1u
M34 net0283 SI VDD VDD PMOS w=6u l=1u
M35 net0283 SE VDD VDD PMOS w=6u l=1u
M38 net0275 net0283 VDD VDD PMOS w=6u l=1u
M26 Q net66 VDD VDD PMOS w=6u l=1u
M24 net66 net92 VDD VDD PMOS w=6u l=1u
M18 net78 net116 N003 VDD PMOS w=6u l=1u
M17 net78 net74 N004 VDD PMOS w=6u l=1u
M16 N003 net104 VDD VDD PMOS w=6u l=1u
M15 N004 net92 VDD VDD PMOS w=6u l=1u
M14 net92 net78 VDD VDD PMOS w=6u l=1u
M13 net104 net114 VDD VDD PMOS w=6u l=1u
M12 N002 net104 VDD VDD PMOS w=6u l=1u
M11 N001 net0275 VDD VDD PMOS w=6u l=1u
M10 net114 net116 N002 VDD PMOS w=6u l=1u
M9 net114 net74 N001 VDD PMOS w=6u l=1u
M8 net116 net74 VDD VDD PMOS w=6u l=1u
M7 net74 CK VDD VDD PMOS w=6u l=1u
M41 N010 net0283 VSS VSS NMOS w=2u l=1u
M40 net0275 net0287 N010 VSS NMOS w=2u l=1u
M29 net0367 SE VSS VSS NMOS w=2u l=1u
M30 N011 net0367 VSS VSS NMOS w=2u l=1u
M31 net0287 D N011 VSS NMOS w=2u l=1u
M36 net0283 SE N005 VSS NMOS w=2u l=1u
M37 N005 SI VSS VSS NMOS w=2u l=1u
M27 Q net66 VSS VSS NMOS w=2u l=1u
M25 net66 net92 VSS VSS NMOS w=2u l=1u
M23 net78 net74 N008 VSS NMOS w=2u l=1u
M22 N008 net104 VSS VSS NMOS w=2u l=1u
M21 net78 net116 N009 VSS NMOS w=2u l=1u
M20 N009 net92 VSS VSS NMOS w=2u l=1u
M19 net92 net78 VSS VSS NMOS w=2u l=1u
M6 net116 net74 VSS VSS NMOS w=2u l=1u
M5 net74 CK VSS VSS NMOS w=2u l=1u
M4 net104 net114 VSS VSS NMOS w=2u l=1u
M3 N007 net104 VSS VSS NMOS w=2u l=1u
M2 net114 net74 N007 VSS NMOS w=2u l=1u
M1 N006 net0275 VSS VSS NMOS w=2u l=1u
M0 net114 net116 N006 VSS NMOS w=2u l=1u
.ends sdff1

.subckt sff1 CK D Q S VDD VSS
M28 net104 S VDD VDD PMOS w=6u l=1u
M31 net92 S VDD VDD PMOS w=6u l=1u
M26 Q net66 VDD VDD PMOS w=6u l=1u
M24 net66 net92 VDD VDD PMOS w=6u l=1u
M18 net78 net116 N003 VDD PMOS w=6u l=1u
M17 net78 net74 N004 VDD PMOS w=6u l=1u
M16 N003 net104 VDD VDD PMOS w=6u l=1u
M15 N004 net92 VDD VDD PMOS w=6u l=1u
M14 net92 net78 VDD VDD PMOS w=6u l=1u
M13 net104 net114 VDD VDD PMOS w=6u l=1u
M12 N002 net104 VDD VDD PMOS w=6u l=1u
M11 N001 D VDD VDD PMOS w=6u l=1u
M10 net114 net116 N002 VDD PMOS w=6u l=1u
M9 net114 net74 N001 VDD PMOS w=6u l=1u
M8 net116 net74 VDD VDD PMOS w=6u l=1u
M7 net74 CK VDD VDD PMOS w=6u l=1u
M27 Q net66 VSS VSS NMOS w=2u l=1u
M25 net66 net92 VSS VSS NMOS w=2u l=1u
M30 N010 net78 VSS VSS NMOS w=2u l=1u
M23 net78 net74 N008 VSS NMOS w=2u l=1u
M22 N008 net104 VSS VSS NMOS w=2u l=1u
M21 net78 net116 N009 VSS NMOS w=2u l=1u
M20 N009 net92 VSS VSS NMOS w=2u l=1u
M19 net92 S N010 VSS NMOS w=2u l=1u
M29 N007 net114 VSS VSS NMOS w=2u l=1u
M6 net116 net74 VSS VSS NMOS w=2u l=1u
M5 net74 CK VSS VSS NMOS w=2u l=1u
M4 net104 S N007 VSS NMOS w=2u l=1u
M3 N006 net104 VSS VSS NMOS w=2u l=1u
M2 net114 net74 N006 VSS NMOS w=2u l=1u
M1 N005 D VSS VSS NMOS w=2u l=1u
M0 net114 net116 N005 VSS NMOS w=2u l=1u
.ends sff1

.subckt srff1 CK D Q R SE SI VDD VSS
M38 net0184 net0176 VDD VDD PMOS w=6u l=1u
M35 net0176 SE VDD VDD PMOS w=6u l=1u
M34 net0176 SI VDD VDD PMOS w=6u l=1u
M33 net0172 net0268 VDD VDD PMOS w=6u l=1u
M36 net0172 D VDD VDD PMOS w=6u l=1u
M29 net104 R N003 VDD PMOS w=6u l=1u
M31 net92 R N006 VDD PMOS w=6u l=1u
M26 Q net66 VDD VDD PMOS w=6u l=1u
M24 net66 net92 VDD VDD PMOS w=6u l=1u
M18 net78 net116 N004 VDD PMOS w=6u l=1u
M17 net78 net74 N005 VDD PMOS w=6u l=1u
M16 N004 net104 VDD VDD PMOS w=6u l=1u
M15 N005 net92 VDD VDD PMOS w=6u l=1u
M14 N006 net78 VDD VDD PMOS w=6u l=1u
M13 N003 net114 VDD VDD PMOS w=6u l=1u
M12 N002 net104 VDD VDD PMOS w=6u l=1u
M11 N001 net0184 VDD VDD PMOS w=6u l=1u
M10 net114 net116 N002 VDD PMOS w=6u l=1u
M9 net114 net74 N001 VDD PMOS w=6u l=1u
M8 net116 net74 VDD VDD PMOS w=6u l=1u
M7 net74 CK VDD VDD PMOS w=6u l=1u
M39 net0184 net0172 VDD VDD PMOS w=6u l=1u
M32 net0268 SE VDD VDD PMOS w=6u l=1u
M37 net0172 D N013 VSS NMOS w=2u l=1u
M40 N013 net0268 VSS VSS NMOS w=2u l=1u
M41 N007 SI VSS VSS NMOS w=2u l=1u
M42 net0176 SE N007 VSS NMOS w=2u l=1u
M43 net0268 SE VSS VSS NMOS w=2u l=1u
M44 N008 net0176 VSS VSS NMOS w=2u l=1u
M45 net0184 net0172 N008 VSS NMOS w=2u l=1u
M27 Q net66 VSS VSS NMOS w=2u l=1u
M25 net66 net92 VSS VSS NMOS w=2u l=1u
M23 net78 net74 N011 VSS NMOS w=2u l=1u
M22 N011 net104 VSS VSS NMOS w=2u l=1u
M21 net78 net116 N012 VSS NMOS w=2u l=1u
M20 N012 net92 VSS VSS NMOS w=2u l=1u
M19 net92 net78 VSS VSS NMOS w=2u l=1u
M30 net92 R VSS VSS NMOS w=2u l=1u
M28 net104 R VSS VSS NMOS w=2u l=1u
M6 net116 net74 VSS VSS NMOS w=2u l=1u
M5 net74 CK VSS VSS NMOS w=2u l=1u
M4 net104 net114 VSS VSS NMOS w=2u l=1u
M3 N010 net104 VSS VSS NMOS w=2u l=1u
M2 net114 net74 N010 VSS NMOS w=2u l=1u
M1 N009 net0184 VSS VSS NMOS w=2u l=1u
M0 net114 net116 N009 VSS NMOS w=2u l=1u
.ends srff1

.subckt ssff1 CK D Q S SE SI VDD VSS
M33 net0178 D VDD VDD PMOS w=6u l=1u
M34 net0178 net0274 VDD VDD PMOS w=6u l=1u
M35 net0174 SI VDD VDD PMOS w=6u l=1u
M36 net0174 SE VDD VDD PMOS w=6u l=1u
M38 net0166 net0174 VDD VDD PMOS w=6u l=1u
M28 net104 S VDD VDD PMOS w=6u l=1u
M31 net92 S VDD VDD PMOS w=6u l=1u
M26 Q net66 VDD VDD PMOS w=6u l=1u
M24 net66 net92 VDD VDD PMOS w=6u l=1u
M18 net78 net116 N003 VDD PMOS w=6u l=1u
M17 net78 net74 N004 VDD PMOS w=6u l=1u
M16 N003 net104 VDD VDD PMOS w=6u l=1u
M15 N004 net92 VDD VDD PMOS w=6u l=1u
M14 net92 net78 VDD VDD PMOS w=6u l=1u
M13 net104 net114 VDD VDD PMOS w=6u l=1u
M12 N002 net104 VDD VDD PMOS w=6u l=1u
M11 N001 net0166 VDD VDD PMOS w=6u l=1u
M10 net114 net116 N002 VDD PMOS w=6u l=1u
M9 net114 net74 N001 VDD PMOS w=6u l=1u
M8 net116 net74 VDD VDD PMOS w=6u l=1u
M7 net74 CK VDD VDD PMOS w=6u l=1u
M32 net0274 SE VDD VDD PMOS w=6u l=1u
M39 net0166 net0178 VDD VDD PMOS w=6u l=1u
M41 N006 net0174 VSS VSS NMOS w=2u l=1u
M40 net0166 net0178 N006 VSS NMOS w=2u l=1u
M37 net0274 SE VSS VSS NMOS w=2u l=1u
M42 N013 net0274 VSS VSS NMOS w=2u l=1u
M43 net0178 D N013 VSS NMOS w=2u l=1u
M44 net0174 SE N005 VSS NMOS w=2u l=1u
M45 N005 SI VSS VSS NMOS w=2u l=1u
M27 Q net66 VSS VSS NMOS w=2u l=1u
M25 net66 net92 VSS VSS NMOS w=2u l=1u
M30 N012 net78 VSS VSS NMOS w=2u l=1u
M23 net78 net74 N010 VSS NMOS w=2u l=1u
M22 N010 net104 VSS VSS NMOS w=2u l=1u
M21 net78 net116 N011 VSS NMOS w=2u l=1u
M20 N011 net92 VSS VSS NMOS w=2u l=1u
M19 net92 S N012 VSS NMOS w=2u l=1u
M29 N009 net114 VSS VSS NMOS w=2u l=1u
M6 net116 net74 VSS VSS NMOS w=2u l=1u
M5 net74 CK VSS VSS NMOS w=2u l=1u
M4 net104 S N009 VSS NMOS w=2u l=1u
M3 N008 net104 VSS VSS NMOS w=2u l=1u
M2 net114 net74 N008 VSS NMOS w=2u l=1u
M1 N007 net0166 VSS VSS NMOS w=2u l=1u
M0 net114 net116 N007 VSS NMOS w=2u l=1u
.ends ssff1
